module bcd7seg(
  input  [3:0] b,               // 输入4位二进制
  output reg [7:0] h            // 输出7段数码管信号
);
  always @(*) begin
    case (b)
        4'b0000: h = 8'b00000011;  // 0
        4'b0001: h = 8'b10011111;  // 1
        4'b0010: h = 8'b00100101;  // 2
        4'b0011: h = 8'b00001101;  // 3
        4'b0100: h = 8'b10011001;  // 4
        4'b0101: h = 8'b01001001;  // 5
        4'b0110: h = 8'b01000001;  // 6
        4'b0111: h = 8'b00011111;  // 7
        4'b1000: h = 8'b00000001;  // 8
        4'b1001: h = 8'b00001001;  // 9
        4'b1010: h = 8'b00010001;  // A
        4'b1011: h = 8'b11000001;  // B
        4'b1100: h = 8'b01100011;  // C
        4'b1101: h = 8'b10000101;  // D
        4'b1110: h = 8'b01100001;  // E
        4'b1111: h = 8'b01110001;  // F
        default: h = 8'b11111111;  // 默认显示空白
    endcase
  end
endmodule
